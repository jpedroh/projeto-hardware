module CPU (clock, reset);

input clock;
input reset;

endmodule