
        {
            "id": "814631019994546216",
            "name": "Chefia da FIR Amazônica",
        },
        {
            "id": "814631152564174888",
            "name": "Chefia da FIR Recife",
        },
        {
            "id": "814631180489064499",
            "name": "Chefia da FIR Curitiba",
        },
        {
            "id": "814631202186723438",
            "name": "Chefia da FIR Brasília",
        },
        {
            "id": "814631220633403402",
            "name": "Chefia da FIR Atlântico",
        },
        {
            "id": "814631238614777868",
            "name": "Chefia do SRPV São Paulo",
        }